
`timescale 1ns / 1ps
//*************************************************************************
//   > 文件名: inst_rom.v
//   > 描述  ：异步指令存储器模块，采用寄存器搭建而成，类似寄存器堆
//   >         内嵌好指令，只读，异步读
//   > 作者  : LOONGSON
//   > 日期  : 2016-04-14
//*************************************************************************
module inst_rom(
    input      [4 :0] addr, // 指令地址
    output reg [31:0] inst       // 指令
  );

  wire [31:0] inst_rom[19:0];  // 指令存储器，字节地址7'b000_0000~7'b111_1111
  //------------- 指令编码 ---------|指令地址|--- 汇编指令 -----|- 指令结果 -----//
  assign inst_rom[ 0] = 32'h24010001; // 00H: addiu $1 ,$0,#1   | $1 = 0000_0001H
  assign inst_rom[ 1] = 32'h00011100; // 04H: sll   $2 ,$1,#4   | $2 = 0000_0010H
  assign inst_rom[ 2] = 32'h00411821; // 08H: addu  $3 ,$2,$1   | $3 = 0000_0011H
  assign inst_rom[ 3] = 32'h00022082; // 0CH: srl   $4 ,$2,#2   | $4 = 0000_0004H
  assign inst_rom[ 4] = 32'h00642823; // 10H: subu  $5 ,$3,$4   | $5 = 0000_000DH
  assign inst_rom[ 5] = 32'hAC250013; // 14H: sw    $5 ,#19($1) | Mem[0000_0014H] = 0000_000DH
  assign inst_rom[ 6] = 32'h00A23027; // 18H: nor   $6 ,$5,$2   | $6 = FFFF_FFE2H
  assign inst_rom[ 7] = 32'h00C33825; // 1CH: or    $7 ,$6,$3   | $7 = FFFF_FFF3H
  assign inst_rom[ 8] = 32'h00E64026; // 20H: xor   $8 ,$7,$6   | $8 = 0000_0011H
  assign inst_rom[ 9] = 32'hAC08001C; // 24H: sw    $8 ,#28($0) | Mem[0000_001CH] = 0000_0011H
  assign inst_rom[10] = 32'h00C7482A; // 28H: slt   $9 ,$6,$7   | $9 = 0000_0001H
  assign inst_rom[11] = 32'h11210002; // 2CH: beq   $9 ,$1,#2   | 跳转到指令34H
  assign inst_rom[12] = 32'h24010004; // 30H: addiu $1 ,$0,#4   | 不执行
  assign inst_rom[13] = 32'h8C2A0013; // 34H: lw    $10,#19($1) | $10 = 0000_000DH
  assign inst_rom[14] = 32'h15450003; // 38H: bne   $10,$5,#3   | 不跳转
  assign inst_rom[15] = 32'h00415824; // 3CH: and   $11,$2,$1   | $11 = 0000_0000H
  assign inst_rom[16] = 32'hAC0B001C; // 40H: sw    $11,#28($0) | Men[0000_001CH] = 0000_0000H
  assign inst_rom[17] = 32'hAC040010; // 44H: sw    $4 ,#16($0) | Mem[0000_0010H] = 0000_0004H
  assign inst_rom[18] = 32'h3C0C000C; // 48H: lui   $12,#12     | [R12] = 000C_0000H
  assign inst_rom[19] = 32'h08000000; // 4CH: j     00H         | 跳转指令00H

  //读指令,取4字节
  always @(*) begin
    case (addr)
      5'd0 :
        inst <= inst_rom[0 ];
      5'd1 :
        inst <= inst_rom[1 ];
      5'd2 :
        inst <= inst_rom[2 ];
      5'd3 :
        inst <= inst_rom[3 ];
      5'd4 :
        inst <= inst_rom[4 ];
      5'd5 :
        inst <= inst_rom[5 ];
      5'd6 :
        inst <= inst_rom[6 ];
      5'd7 :
        inst <= inst_rom[7 ];
      5'd8 :
        inst <= inst_rom[8 ];
      5'd9 :
        inst <= inst_rom[9 ];
      5'd10:
        inst <= inst_rom[10];
      5'd11:
        inst <= inst_rom[11];
      5'd12:
        inst <= inst_rom[12];
      5'd13:
        inst <= inst_rom[13];
      5'd14:
        inst <= inst_rom[14];
      5'd15:
        inst <= inst_rom[15];
      5'd16:
        inst <= inst_rom[16];
      5'd17:
        inst <= inst_rom[17];
      5'd18:
        inst <= inst_rom[18];
      5'd19:
        inst <= inst_rom[19];
      default:
        inst <= 32'd0;
    endcase
  end
endmodule
